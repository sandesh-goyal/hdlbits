module top_module (
    input a, b, c, d, e,
    output [24:0] out );//

    // The output is XNOR of two vectors created by 
    // concatenating and replicating the five inputs.
    // assign out = ~{ ... } ^ { ... };
    wire [24:0] out1, out3;
    wire [4:0] out2;
    assign out1 = {{5{a}}, {5{b}}, {5{c}}, {5{d}}, {5{e}}};
    assign out2 = {a,b,c,d,e};
    assign out3 = {5{a,b,c,d,e}};
    assign out = ~(out1 ^ out3);

endmodule
